/**
 * pll.v
 * PLL configuration
 * This Verilog module was generated automatically using the icepll tool from the IceStorm project.
 */

module pll(
    input  clk_in,
    output clk_out,
    output locked
    );

SB_PLL40_CORE #(
        .FEEDBACK_PATH("SIMPLE"),
        .DIVR(4'b0000),        // DIVR =  0
        .DIVF(7'b1001111),     // DIVF = 79
        .DIVQ(3'b100),         // DIVQ =  4
        .FILTER_RANGE(3'b001)  // FILTER_RANGE = 1
    ) uut (
        .LOCK(locked),
        .RESETB(1'b1),
        .BYPASS(1'b0),
        .REFERENCECLK(clk_in),
        .PLLOUTCORE(clk_out)
        );

endmodule
